`timescale 1ps/1ps
`default_nettype none

module axi_crossbar_top#(
    parameter AXI_ID_W   = 4,
    parameter AXI_DATA_W = 32,
    parameter AXI_ADDR_W = 32,

    parameter MST_NB     = 3,
    parameter SLV_NB     = 3,

    parameter MST_PIPELINE = 1,
    parameter SLV_PIPELINE = 1,

    //Master0 Configuration
    parameter MST0_OSTDREQ_NUM = 4,
    parameter MST0_OSTDREQ_SIZE = 1,
    parameter MST0_PRIORITY = 0,
    parameter [SLV_NB-1:0] MST0_ROUTES = 3'b1_1_1,
    parameter [AXI_ID_W-1:0] MST0_ID_MASK = 4'b01_00,

    //Master1 Configuration
    parameter MST1_OSTDREQ_NUM = 4,
    parameter MST1_OSTDREQ_SIZE = 1,
    parameter MST1_PRIORITY = 0,
    parameter [SLV_NB-1:0] MST1_ROUTES = 3'b1_1_1,
    parameter [AXI_ID_W-1:0] MST1_ID_MASK = 4'b10_00,

    //Master2 Configuration
    parameter MST2_OSTDREQ_NUM = 4,
    parameter MST2_OSTDREQ_SIZE = 1,
    parameter MST2_PRIORITY = 0,
    parameter [SLV_NB-1:0] MST2_ROUTES = 3'b1_1_1,
    parameter [AXI_ID_W-1:0] MST2_ID_MASK = 4'b11_00,

    //SLV0 Configuration
    parameter SLV0_START_ADDR = 0,
    parameter SLV0_END_ADDR = 4095,
    parameter SLV0_OSTDREQ_NUM = 4,
    parameter SLV0_OSTDREQ_SIZE = 1,
    parameter SLV0_PRIORITY = 0,

    //SLV1 Configuration
    parameter SLV1_START_ADDR = 4096,
    parameter SLV1_END_ADDR = 8191,
    parameter SLV1_OSTDREQ_NUM = 4,
    parameter SLV1_OSTDREQ_SIZE = 1,
    parameter SLV1_PRIORITY = 0,

    //SLV2 Configuration
    parameter SLV2_START_ADDR = 8192,
    parameter SLV2_END_ADDR = 12287,
    parameter SLV2_OSTDREQ_NUM = 4,
    parameter SLV2_OSTDREQ_SIZE = 1,
    parameter SLV2_PRIORITY = 0,

    // Channels' width (concatenated)
    parameter AWCH_W = 49,
    parameter WCH_W  = 43,
    parameter BCH_W  = 8,
    parameter ARCH_W = 49,
    parameter RCH_W  = 41,    
    
    //CAM parameters
    parameter CAM_ADDR_WIDTH = 4    
    )(
    //crossbar inner signal
    input  wire                       aclk,
    input  wire                       aresetn,
    input  wire                       srst,

    //mst0 interface
    input  wire                       mst0_aclk,
    input  wire                       mst0_aresetn,
    input  wire                       mst0_srst,
    input  wire                       mst0_awvalid,
    output logic                      mst0_awready,
    input  wire  [AXI_ADDR_W    -1:0] mst0_awaddr,
    input  wire  [4             -1:0] mst0_awlen,
    input  wire  [3             -1:0] mst0_awsize,
    input  wire  [2             -1:0] mst0_awburst,
    input  wire  [2             -1:0] mst0_awlock,
    input  wire  [AXI_ID_W      -1:0] mst0_awid,
    input  wire                       mst0_wvalid,
    output logic                      mst0_wready,
    input  wire                       mst0_wlast,
    input  wire  [AXI_DATA_W    -1:0] mst0_wdata,
    input  wire  [AXI_DATA_W/8  -1:0] mst0_wstrb,
    input  wire  [AXI_ID_W      -1:0] mst0_wid,
    output logic                      mst0_bvalid,
    input  wire                       mst0_bready,
    output logic [AXI_ID_W      -1:0] mst0_bid,
    output logic [2             -1:0] mst0_bresp,
    input  wire                       mst0_arvalid,
    output logic                      mst0_arready,
    input  wire  [AXI_ADDR_W    -1:0] mst0_araddr,
    input  wire  [4             -1:0] mst0_arlen,
    input  wire  [3             -1:0] mst0_arsize,
    input  wire  [2             -1:0] mst0_arburst,
    input  wire  [2             -1:0] mst0_arlock,
    input  wire  [AXI_ID_W      -1:0] mst0_arid,
    output logic                      mst0_rvalid,
    input  wire                       mst0_rready,
    output logic [AXI_ID_W      -1:0] mst0_rid,
    output logic [2             -1:0] mst0_rresp,
    output logic [AXI_DATA_W    -1:0] mst0_rdata,
    output logic                      mst0_rlast,

    //mst1 interface
    input  wire                       mst1_aclk,
    input  wire                       mst1_aresetn,
    input  wire                       mst1_srst,
    input  wire                       mst1_awvalid,
    output logic                      mst1_awready,
    input  wire  [AXI_ADDR_W    -1:0] mst1_awaddr,
    input  wire  [4             -1:0] mst1_awlen,
    input  wire  [3             -1:0] mst1_awsize,
    input  wire  [2             -1:0] mst1_awburst,
    input  wire  [2             -1:0] mst1_awlock,
    input  wire  [AXI_ID_W      -1:0] mst1_awid,
    input  wire                       mst1_wvalid,
    output logic                      mst1_wready,
    input  wire                       mst1_wlast,
    input  wire  [AXI_DATA_W    -1:0] mst1_wdata,
    input  wire  [AXI_DATA_W/8  -1:0] mst1_wstrb,
    input  wire  [AXI_ID_W      -1:0] mst1_wid,
    output logic                      mst1_bvalid,
    input  wire                       mst1_bready,
    output logic [AXI_ID_W      -1:0] mst1_bid,
    output logic [2             -1:0] mst1_bresp,
    input  wire                       mst1_arvalid,
    output logic                      mst1_arready,
    input  wire  [AXI_ADDR_W    -1:0] mst1_araddr,
    input  wire  [4             -1:0] mst1_arlen,
    input  wire  [3             -1:0] mst1_arsize,
    input  wire  [2             -1:0] mst1_arburst,
    input  wire  [2             -1:0] mst1_arlock,
    input  wire  [AXI_ID_W      -1:0] mst1_arid,
    output logic                      mst1_rvalid,
    input  wire                       mst1_rready,
    output logic [AXI_ID_W      -1:0] mst1_rid,
    output logic [2             -1:0] mst1_rresp,
    output logic [AXI_DATA_W    -1:0] mst1_rdata,
    output logic                      mst1_rlast,

    //mst2 interface
    input  wire                       mst2_aclk,
    input  wire                       mst2_aresetn,
    input  wire                       mst2_srst,
    input  wire                       mst2_awvalid,
    output logic                      mst2_awready,
    input  wire  [AXI_ADDR_W    -1:0] mst2_awaddr,
    input  wire  [4             -1:0] mst2_awlen,
    input  wire  [3             -1:0] mst2_awsize,
    input  wire  [2             -1:0] mst2_awburst,
    input  wire  [2             -1:0] mst2_awlock,
    input  wire  [AXI_ID_W      -1:0] mst2_awid,
    input  wire                       mst2_wvalid,
    output logic                      mst2_wready,
    input  wire                       mst2_wlast,
    input  wire  [AXI_DATA_W    -1:0] mst2_wdata,
    input  wire  [AXI_DATA_W/8  -1:0] mst2_wstrb,
    input  wire  [AXI_ID_W      -1:0] mst2_wid,
    output logic                      mst2_bvalid,
    input  wire                       mst2_bready,
    output logic [AXI_ID_W      -1:0] mst2_bid,
    output logic [2             -1:0] mst2_bresp,
    input  wire                       mst2_arvalid,
    output logic                      mst2_arready,
    input  wire  [AXI_ADDR_W    -1:0] mst2_araddr,
    input  wire  [4             -1:0] mst2_arlen,
    input  wire  [3             -1:0] mst2_arsize,
    input  wire  [2             -1:0] mst2_arburst,
    input  wire  [2             -1:0] mst2_arlock,
    input  wire  [AXI_ID_W      -1:0] mst2_arid,
    output logic                      mst2_rvalid,
    input  wire                       mst2_rready,
    output logic [AXI_ID_W      -1:0] mst2_rid,
    output logic [2             -1:0] mst2_rresp,
    output logic [AXI_DATA_W    -1:0] mst2_rdata,
    output logic                      mst2_rlast,

    //slv0 interface
    input  wire                       slv0_aclk,
    input  wire                       slv0_aresetn,
    input  wire                       slv0_srst,
    output logic                      slv0_awvalid,
    input  wire                       slv0_awready,
    output logic [AXI_ADDR_W    -1:0] slv0_awaddr,
    output logic [4             -1:0] slv0_awlen,
    output logic [3             -1:0] slv0_awsize,
    output logic [2             -1:0] slv0_awburst,
    output logic [2             -1:0] slv0_awlock,
    output logic [AXI_ID_W      -1:0] slv0_awid,
    output logic                      slv0_wvalid,
    input  wire                       slv0_wready,
    output logic                      slv0_wlast,
    output logic [AXI_DATA_W    -1:0] slv0_wdata,
    output logic [AXI_DATA_W/8  -1:0] slv0_wstrb,
    output logic [AXI_ID_W      -1:0] slv0_wid,
    input  wire                       slv0_bvalid,
    output logic                      slv0_bready,
    input  wire  [AXI_ID_W      -1:0] slv0_bid,
    input  wire  [2             -1:0] slv0_bresp,
    output logic                      slv0_arvalid,
    input  wire                       slv0_arready,
    output logic [AXI_ADDR_W    -1:0] slv0_araddr,
    output logic [4             -1:0] slv0_arlen,
    output logic [3             -1:0] slv0_arsize,
    output logic [2             -1:0] slv0_arburst,
    output logic [2             -1:0] slv0_arlock,
    output logic [AXI_ID_W      -1:0] slv0_arid,
    input  wire                       slv0_rvalid,
    output logic                      slv0_rready,
    input  wire  [AXI_ID_W      -1:0] slv0_rid,
    input  wire  [2             -1:0] slv0_rresp,
    input  wire  [AXI_DATA_W    -1:0] slv0_rdata,
    input  wire                       slv0_rlast,

    //slv1 interface
    input  wire                       slv1_aclk,
    input  wire                       slv1_aresetn,
    input  wire                       slv1_srst,
    output logic                      slv1_awvalid,
    input  wire                       slv1_awready,
    output logic [AXI_ADDR_W    -1:0] slv1_awaddr,
    output logic [4             -1:0] slv1_awlen,
    output logic [3             -1:0] slv1_awsize,
    output logic [2             -1:0] slv1_awburst,
    output logic [2             -1:0] slv1_awlock,
    output logic [AXI_ID_W      -1:0] slv1_awid,
    output logic                      slv1_wvalid,
    input  wire                       slv1_wready,
    output logic                      slv1_wlast,
    output logic [AXI_DATA_W    -1:0] slv1_wdata,
    output logic [AXI_DATA_W/8  -1:0] slv1_wstrb,
    output logic [AXI_ID_W      -1:0] slv1_wid,
    input  wire                       slv1_bvalid,
    output logic                      slv1_bready,
    input  wire  [AXI_ID_W      -1:0] slv1_bid,
    input  wire  [2             -1:0] slv1_bresp,
    output logic                      slv1_arvalid,
    input  wire                       slv1_arready,
    output logic [AXI_ADDR_W    -1:0] slv1_araddr,
    output logic [4             -1:0] slv1_arlen,
    output logic [3             -1:0] slv1_arsize,
    output logic [2             -1:0] slv1_arburst,
    output logic [2             -1:0] slv1_arlock,
    output logic [AXI_ID_W      -1:0] slv1_arid,
    input  wire                       slv1_rvalid,
    output logic                      slv1_rready,
    input  wire  [AXI_ID_W      -1:0] slv1_rid,
    input  wire  [2             -1:0] slv1_rresp,
    input  wire  [AXI_DATA_W    -1:0] slv1_rdata,
    input  wire                       slv1_rlast,

    //slv2 interface
    input  wire                       slv2_aclk,
    input  wire                       slv2_aresetn,
    input  wire                       slv2_srst,
    output logic                      slv2_awvalid,
    input  wire                       slv2_awready,
    output logic [AXI_ADDR_W    -1:0] slv2_awaddr,
    output logic [4             -1:0] slv2_awlen,
    output logic [3             -1:0] slv2_awsize,
    output logic [2             -1:0] slv2_awburst,
    output logic [2             -1:0] slv2_awlock,
    output logic [AXI_ID_W      -1:0] slv2_awid,
    output logic                      slv2_wvalid,
    input  wire                       slv2_wready,
    output logic                      slv2_wlast,
    output logic [AXI_DATA_W    -1:0] slv2_wdata,
    output logic [AXI_DATA_W/8  -1:0] slv2_wstrb,
    output logic [AXI_ID_W      -1:0] slv2_wid,
    input  wire                       slv2_bvalid,
    output logic                      slv2_bready,
    input  wire  [AXI_ID_W      -1:0] slv2_bid,
    input  wire  [2             -1:0] slv2_bresp,
    output logic                      slv2_arvalid,
    input  wire                       slv2_arready,
    output logic [AXI_ADDR_W    -1:0] slv2_araddr,
    output logic [4             -1:0] slv2_arlen,
    output logic [3             -1:0] slv2_arsize,
    output logic [2             -1:0] slv2_arburst,
    output logic [2             -1:0] slv2_arlock,
    output logic [AXI_ID_W      -1:0] slv2_arid,
    input  wire                       slv2_rvalid,
    output logic                      slv2_rready,
    input  wire  [AXI_ID_W      -1:0] slv2_rid,
    input  wire  [2             -1:0] slv2_rresp,
    input  wire  [AXI_DATA_W    -1:0] slv2_rdata,
    input  wire                       slv2_rlast    
    );
    //local declaration
    localparam MST_ROUTES = {MST2_ROUTES,
                             MST1_ROUTES,
                             MST0_ROUTES};

    logic [MST_NB            -1:0] i_awvalid;
    logic [MST_NB            -1:0] i_awready;
    logic [MST_NB*AWCH_W     -1:0] i_awch;
    logic [MST_NB            -1:0] i_wvalid;
    logic [MST_NB            -1:0] i_wready;
    logic [MST_NB            -1:0] i_wlast;
    logic [MST_NB*WCH_W      -1:0] i_wch;
    logic [MST_NB            -1:0] i_bvalid;
    logic [MST_NB            -1:0] i_bready;
    logic [MST_NB*BCH_W      -1:0] i_bch;
    logic [MST_NB            -1:0] i_arvalid;
    logic [MST_NB            -1:0] i_arready;
    logic [MST_NB*ARCH_W     -1:0] i_arch;
    logic [MST_NB            -1:0] i_rvalid;
    logic [MST_NB            -1:0] i_rready;
    logic [MST_NB            -1:0] i_rlast;
    logic [MST_NB*RCH_W      -1:0] i_rch;
    logic [SLV_NB            -1:0] o_awvalid;
    logic [SLV_NB            -1:0] o_awready;
    logic [SLV_NB*AWCH_W     -1:0] o_awch;
    logic [SLV_NB            -1:0] o_wvalid;
    logic [SLV_NB            -1:0] o_wready;
    logic [SLV_NB            -1:0] o_wlast;
    logic [SLV_NB*WCH_W      -1:0] o_wch;
    logic [SLV_NB            -1:0] o_bvalid;
    logic [SLV_NB            -1:0] o_bready;
    logic [SLV_NB*BCH_W      -1:0] o_bch;
    logic [SLV_NB            -1:0] o_arvalid;
    logic [SLV_NB            -1:0] o_arready;
    logic [SLV_NB*ARCH_W     -1:0] o_arch;
    logic [SLV_NB            -1:0] o_rvalid;
    logic [SLV_NB            -1:0] o_rready;
    logic [SLV_NB            -1:0] o_rlast;
    logic [SLV_NB*RCH_W      -1:0] o_rch;           

    ////////////////////////////////
    //mst0 interface
    ///////////////////////////////
    axi_crossbar_mst_if #(
        .AXI_ADDR_W        (AXI_ADDR_W),
        .AXI_ID_W          (AXI_ID_W),
        .AXI_DATA_W        (AXI_DATA_W),
        .MST_OSTDREQ_NUM   (MST0_OSTDREQ_NUM),
        .MST_OSTDREQ_SIZE  (MST0_OSTDREQ_SIZE),
        .AWCH_W            (AWCH_W),
        .WCH_W             (WCH_W),
        .BCH_W             (BCH_W),
        .ARCH_W            (ARCH_W),
        .RCH_W             (RCH_W),
        .MST_ID_MASK       (MST0_ID_MASK)
    )
        mst0_if(
        .i_aclk       (mst0_aclk),
        .i_aresetn    (mst0_aresetn),
        .i_srst       (mst0_srst),
        //interface from mst
        .i_awvalid    (mst0_awvalid),
        .i_awready    (mst0_awready),
        .i_awaddr     (mst0_awaddr),
        .i_awlen      (mst0_awlen),
        .i_awsize     (mst0_awsize),
        .i_awburst    (mst0_awburst),
        .i_awlock     (mst0_awlock),
        .i_awid       (mst0_awid),
        .i_wvalid     (mst0_wvalid),
        .i_wready     (mst0_wready),
        .i_wlast      (mst0_wlast ),
        .i_wid        (mst0_wid),
        .i_wdata      (mst0_wdata),
        .i_wstrb      (mst0_wstrb),
        .i_bvalid     (mst0_bvalid),
        .i_bready     (mst0_bready),
        .i_bid        (mst0_bid),
        .i_bresp      (mst0_bresp),
        .i_arvalid    (mst0_arvalid),
        .i_arready    (mst0_arready),
        .i_araddr     (mst0_araddr),
        .i_arlen      (mst0_arlen),
        .i_arsize     (mst0_arsize),
        .i_arburst    (mst0_arburst),
        .i_arlock     (mst0_arlock),
        .i_arid       (mst0_arid),
        .i_rvalid     (mst0_rvalid),
        .i_rready     (mst0_rready),
        .i_rid        (mst0_rid),
        .i_rresp      (mst0_rresp),
        .i_rdata      (mst0_rdata),
        .i_rlast      (mst0_rlast),
        //interface to axi switch
        .o_aclk       (aclk),
        .o_aresetn    (aresetn),
        .o_srst       (srst),
        .o_awvalid    (i_awvalid[0]),
        .o_awready    (i_awready[0]),
        .o_awch       (i_awch[0*AWCH_W+:AWCH_W]),
        .o_wvalid     (i_wvalid[0]),
        .o_wready     (i_wready[0]),
        .o_wlast      (i_wlast[0]),
        .o_wch        (i_wch[0*WCH_W+:WCH_W]),
        .o_bvalid     (i_bvalid[0]),
        .o_bready     (i_bready[0]),
        .o_bch        (i_bch[0*BCH_W+:BCH_W]),
        .o_arvalid    (i_arvalid[0]),
        .o_arready    (i_arready[0]),
        .o_arch       (i_arch[0*ARCH_W+:ARCH_W]),
        .o_rvalid     (i_rvalid[0]),
        .o_rready     (i_rready[0]),
        .o_rlast      (i_rlast[0]),
        .o_rch        (i_rch[0*RCH_W+:RCH_W])
    );

    ////////////////////////////////
    //mst1 interface
    ///////////////////////////////
    axi_crossbar_mst_if #(
        .AXI_ADDR_W        (AXI_ADDR_W),
        .AXI_ID_W          (AXI_ID_W),
        .AXI_DATA_W        (AXI_DATA_W),
        .MST_OSTDREQ_NUM   (MST1_OSTDREQ_NUM),
        .MST_OSTDREQ_SIZE  (MST1_OSTDREQ_SIZE),
        .AWCH_W            (AWCH_W),
        .WCH_W             (WCH_W),
        .BCH_W             (BCH_W),
        .ARCH_W            (ARCH_W),
        .RCH_W             (RCH_W),
        .MST_ID_MASK       (MST1_ID_MASK)
    )
        mst1_if(
        .i_aclk       (mst1_aclk),
        .i_aresetn    (mst1_aresetn),
        .i_srst       (mst1_srst),
        //interface from mst
        .i_awvalid    (mst1_awvalid),
        .i_awready    (mst1_awready),
        .i_awaddr     (mst1_awaddr),
        .i_awlen      (mst1_awlen),
        .i_awsize     (mst1_awsize),
        .i_awburst    (mst1_awburst),
        .i_awlock     (mst1_awlock),
        .i_awid       (mst1_awid),
        .i_wvalid     (mst1_wvalid),
        .i_wready     (mst1_wready),
        .i_wlast      (mst1_wlast ),
        .i_wid        (mst1_wid),
        .i_wdata      (mst1_wdata),
        .i_wstrb      (mst1_wstrb),
        .i_bvalid     (mst1_bvalid),
        .i_bready     (mst1_bready),
        .i_bid        (mst1_bid),
        .i_bresp      (mst1_bresp),
        .i_arvalid    (mst1_arvalid),
        .i_arready    (mst1_arready),
        .i_araddr     (mst1_araddr),
        .i_arlen      (mst1_arlen),
        .i_arsize     (mst1_arsize),
        .i_arburst    (mst1_arburst),
        .i_arlock     (mst1_arlock),
        .i_arid       (mst1_arid),
        .i_rvalid     (mst1_rvalid),
        .i_rready     (mst1_rready),
        .i_rid        (mst1_rid),
        .i_rresp      (mst1_rresp),
        .i_rdata      (mst1_rdata),
        .i_rlast      (mst1_rlast),
        //interface to axi switch
        .o_aclk       (aclk),
        .o_aresetn    (aresetn),
        .o_srst       (srst),
        .o_awvalid    (i_awvalid[1]),
        .o_awready    (i_awready[1]),
        .o_awch       (i_awch[1*AWCH_W+:AWCH_W]),
        .o_wvalid     (i_wvalid[1]),
        .o_wready     (i_wready[1]),
        .o_wlast      (i_wlast[1]),
        .o_wch        (i_wch[1*WCH_W+:WCH_W]),
        .o_bvalid     (i_bvalid[1]),
        .o_bready     (i_bready[1]),
        .o_bch        (i_bch[1*BCH_W+:BCH_W]),
        .o_arvalid    (i_arvalid[1]),
        .o_arready    (i_arready[1]),
        .o_arch       (i_arch[1*ARCH_W+:ARCH_W]),
        .o_rvalid     (i_rvalid[1]),
        .o_rready     (i_rready[1]),
        .o_rlast      (i_rlast[1]),
        .o_rch        (i_rch[1*RCH_W+:RCH_W])
    );

    ////////////////////////////////
    //mst2 interface
    ///////////////////////////////
    axi_crossbar_mst_if #(
        .AXI_ADDR_W        (AXI_ADDR_W),
        .AXI_ID_W          (AXI_ID_W),
        .AXI_DATA_W        (AXI_DATA_W),
        .MST_OSTDREQ_NUM   (MST2_OSTDREQ_NUM),
        .MST_OSTDREQ_SIZE  (MST2_OSTDREQ_SIZE),
        .AWCH_W            (AWCH_W),
        .WCH_W             (WCH_W),
        .BCH_W             (BCH_W),
        .ARCH_W            (ARCH_W),
        .RCH_W             (RCH_W),
        .MST_ID_MASK       (MST2_ID_MASK)
    )
        mst2_if(
        .i_aclk       (mst2_aclk),
        .i_aresetn    (mst2_aresetn),
        .i_srst       (mst2_srst),
        //interface from mst
        .i_awvalid    (mst2_awvalid),
        .i_awready    (mst2_awready),
        .i_awaddr     (mst2_awaddr),
        .i_awlen      (mst2_awlen),
        .i_awsize     (mst2_awsize),
        .i_awburst    (mst2_awburst),
        .i_awlock     (mst2_awlock),
        .i_awid       (mst2_awid),
        .i_wvalid     (mst2_wvalid),
        .i_wready     (mst2_wready),
        .i_wlast      (mst2_wlast ),
        .i_wid        (mst2_wid),
        .i_wdata      (mst2_wdata),
        .i_wstrb      (mst2_wstrb),
        .i_bvalid     (mst2_bvalid),
        .i_bready     (mst2_bready),
        .i_bid        (mst2_bid),
        .i_bresp      (mst2_bresp),
        .i_arvalid    (mst2_arvalid),
        .i_arready    (mst2_arready),
        .i_araddr     (mst2_araddr),
        .i_arlen      (mst2_arlen),
        .i_arsize     (mst2_arsize),
        .i_arburst    (mst2_arburst),
        .i_arlock     (mst2_arlock),
        .i_arid       (mst2_arid),
        .i_rvalid     (mst2_rvalid),
        .i_rready     (mst2_rready),
        .i_rid        (mst2_rid),
        .i_rresp      (mst2_rresp),
        .i_rdata      (mst2_rdata),
        .i_rlast      (mst2_rlast),
        //interface to axi switch
        .o_aclk       (aclk),
        .o_aresetn    (aresetn),
        .o_srst       (srst),
        .o_awvalid    (i_awvalid[2]),
        .o_awready    (i_awready[2]),
        .o_awch       (i_awch[2*AWCH_W+:AWCH_W]),
        .o_wvalid     (i_wvalid[2]),
        .o_wready     (i_wready[2]),
        .o_wlast      (i_wlast[2]),
        .o_wch        (i_wch[2*WCH_W+:WCH_W]),
        .o_bvalid     (i_bvalid[2]),
        .o_bready     (i_bready[2]),
        .o_bch        (i_bch[2*BCH_W+:BCH_W]),
        .o_arvalid    (i_arvalid[2]),
        .o_arready    (i_arready[2]),
        .o_arch       (i_arch[2*ARCH_W+:ARCH_W]),
        .o_rvalid     (i_rvalid[2]),
        .o_rready     (i_rready[2]),
        .o_rlast      (i_rlast[2]),
        .o_rch        (i_rch[2*RCH_W+:RCH_W])
    );    

    ////////////////////////////////
    //switch top
    ///////////////////////////////
    axi_crossbar_switch_top#(
        .AXI_ADDR_W         (AXI_ADDR_W),
        .AXI_ID_W           (AXI_ID_W),
        .AXI_DATA_W         (AXI_DATA_W),
        .MST_NB             (MST_NB),
        .SLV_NB             (SLV_NB),
        .MST_PIPELINE       (MST_PIPELINE),
        .SLV_PIPELINE       (SLV_PIPELINE),
        .MST_ROUTES         (MST_ROUTES),
        .MST_OSTDREQ_NUM    (MST0_OSTDREQ_NUM),
        .MST_OSTDREQ_SIZE   (MST0_OSTDREQ_SIZE),
        .MST0_ID_MASK       (MST0_ID_MASK),
        .MST1_ID_MASK       (MST1_ID_MASK),
        .MST2_ID_MASK       (MST2_ID_MASK),
        .MST0_PRIORITY      (MST0_PRIORITY),
        .MST1_PRIORITY      (MST1_PRIORITY),
        .MST2_PRIORITY      (MST2_PRIORITY),
        .SLV0_PRIORITY      (SLV0_PRIORITY),
        .SLV1_PRIORITY      (SLV1_PRIORITY),
        .SLV2_PRIORITY      (SLV2_PRIORITY),
        .SLV0_START_ADDR    (SLV0_START_ADDR),
        .SLV0_END_ADDR      (SLV0_END_ADDR),
        .SLV1_START_ADDR    (SLV1_START_ADDR),
        .SLV1_END_ADDR      (SLV1_END_ADDR),
        .SLV2_START_ADDR    (SLV2_START_ADDR),
        .SLV2_END_ADDR      (SLV2_END_ADDR),
        .AWCH_W             (AWCH_W),
        .WCH_W              (WCH_W),
        .BCH_W              (BCH_W),
        .ARCH_W             (ARCH_W),
        .RCH_W              (RCH_W),
        .CAM_ADDR_WIDTH     (CAM_ADDR_WIDTH))
    switch_top(
        //axi crossbar inner signal
        .aclk      (aclk),
        .aresetn   (aresetn),
        .srst      (srst),
        //interface from mst interface
        .i_awvalid (i_awvalid),
        .i_awready (i_awready),
        .i_awch    (i_awch),
        .i_wvalid  (i_wvalid),
        .i_wready  (i_wready),
        .i_wlast   (i_wlast),
        .i_wch     (i_wch),
        .i_bvalid  (i_bvalid),
        .i_bready  (i_bready),
        .i_bch     (i_bch),
        .i_arvalid (i_arvalid),
        .i_arready (i_arready),
        .i_arch    (i_arch),
        .i_rvalid  (i_rvalid),
        .i_rready  (i_rready),
        .i_rlast   (i_rlast),
        .i_rch     (i_rch),
        //interface to slv interface
        .o_awvalid (o_awvalid),
        .o_awready (o_awready),
        .o_awch    (o_awch),
        .o_wvalid  (o_wvalid),
        .o_wready  (o_wready),
        .o_wlast   (o_wlast),
        .o_wch     (o_wch),
        .o_bvalid  (o_bvalid),
        .o_bready  (o_bready),
        .o_bch     (o_bch),
        .o_arvalid (o_arvalid),
        .o_arready (o_arready),
        .o_arch    (o_arch),
        .o_rvalid  (o_rvalid),
        .o_rready  (o_rready),
        .o_rlast   (o_rlast),
        .o_rch     (o_rch)
    );

    ////////////////////////////////
    //slv0 interface
    ///////////////////////////////
    axi_crossbar_slv_if#(
        .AXI_ADDR_W       (AXI_ADDR_W),
        .AXI_ID_W         (AXI_ID_W),
        .AXI_DATA_W       (AXI_DATA_W),
        .BASE_ADDR        (SLV0_START_ADDR),
        .SLV_OSTDREQ_NUM  (SLV0_OSTDREQ_NUM),
        .SLV_OSTDREQ_SIZE (SLV0_OSTDREQ_SIZE),
        .AWCH_W           (AWCH_W),
        .WCH_W            (WCH_W),
        .BCH_W            (BCH_W),
        .ARCH_W           (ARCH_W),
        .RCH_W            (RCH_W))
    slv0_if(
         //interface from switch
        .i_aclk       (aclk),
        .i_aresetn    (aresetn),
        .i_srst       (srst),
        .i_awvalid    (o_awvalid[0]),
        .i_awready    (o_awready[0]),
        .i_awch       (o_awch[0*AWCH_W+:AWCH_W]),
        .i_wvalid     (o_wvalid[0]),
        .i_wready     (o_wready[0]),
        .i_wlast      (o_wlast[0]),
        .i_wch        (o_wch[0*WCH_W+:WCH_W]),
        .i_bvalid     (o_bvalid[0]),
        .i_bready     (o_bready[0]),
        .i_bch        (o_bch[0*BCH_W+:BCH_W]),
        .i_arvalid    (o_arvalid[0]),
        .i_arready    (o_arready[0]),
        .i_arch       (o_arch[0*ARCH_W+:ARCH_W]),
        .i_rvalid     (o_rvalid[0]),
        .i_rready     (o_rready[0]),
        .i_rlast      (o_rlast[0]),
        .i_rch        (o_rch[0*RCH_W+:RCH_W]),
        //interface to slave
        .o_aclk       (slv0_aclk),
        .o_aresetn    (slv0_aresetn),
        .o_srst       (slv0_srst),
        .o_awvalid    (slv0_awvalid),
        .o_awready    (slv0_awready),
        .o_awaddr     (slv0_awaddr),
        .o_awlen      (slv0_awlen),
        .o_awsize     (slv0_awsize),
        .o_awburst    (slv0_awburst),
        .o_awlock     (slv0_awlock),
        .o_awid       (slv0_awid),
        .o_wvalid     (slv0_wvalid),
        .o_wready     (slv0_wready),
        .o_wlast      (slv0_wlast),
        .o_wid        (slv0_wid),
        .o_wdata      (slv0_wdata),
        .o_wstrb      (slv0_wstrb),
        .o_bvalid     (slv0_bvalid),
        .o_bready     (slv0_bready),
        .o_bid        (slv0_bid),
        .o_bresp      (slv0_bresp),
        .o_arvalid    (slv0_arvalid),
        .o_arready    (slv0_arready),
        .o_araddr     (slv0_araddr),
        .o_arlen      (slv0_arlen),
        .o_arsize     (slv0_arsize),
        .o_arburst    (slv0_arburst),
        .o_arlock     (slv0_arlock),
        .o_arid       (slv0_arid),
        .o_rvalid     (slv0_rvalid),
        .o_rready     (slv0_rready),
        .o_rid        (slv0_rid),
        .o_rresp      (slv0_rresp),
        .o_rdata      (slv0_rdata),
        .o_rlast      (slv0_rlast)
    );

    ////////////////////////////////
    //slv1 interface
    ///////////////////////////////
    axi_crossbar_slv_if#(
        .AXI_ADDR_W       (AXI_ADDR_W),
        .AXI_ID_W         (AXI_ID_W),
        .AXI_DATA_W       (AXI_DATA_W),
        .BASE_ADDR        (SLV1_START_ADDR),
        .SLV_OSTDREQ_NUM  (SLV1_OSTDREQ_NUM),
        .SLV_OSTDREQ_SIZE (SLV1_OSTDREQ_SIZE),
        .AWCH_W           (AWCH_W),
        .WCH_W            (WCH_W),
        .BCH_W            (BCH_W),
        .ARCH_W           (ARCH_W),
        .RCH_W            (RCH_W)
    )
    slv1_if(
         //interface from switch
        .i_aclk       (aclk),
        .i_aresetn    (aresetn),
        .i_srst       (srst),
        .i_awvalid    (o_awvalid[1]),
        .i_awready    (o_awready[1]),
        .i_awch       (o_awch[1*AWCH_W+:AWCH_W]),
        .i_wvalid     (o_wvalid[1]),
        .i_wready     (o_wready[1]),
        .i_wlast      (o_wlast[1]),
        .i_wch        (o_wch[1*WCH_W+:WCH_W]),
        .i_bvalid     (o_bvalid[1]),
        .i_bready     (o_bready[1]),
        .i_bch        (o_bch[1*BCH_W+:BCH_W]),
        .i_arvalid    (o_arvalid[1]),
        .i_arready    (o_arready[1]),
        .i_arch       (o_arch[1*ARCH_W+:ARCH_W]),
        .i_rvalid     (o_rvalid[1]),
        .i_rready     (o_rready[1]),
        .i_rlast      (o_rlast[1]),
        .i_rch        (o_rch[1*RCH_W+:RCH_W]),
        //interface to slave
        .o_aclk       (slv1_aclk),
        .o_aresetn    (slv1_aresetn),
        .o_srst       (slv1_srst),
        .o_awvalid    (slv1_awvalid),
        .o_awready    (slv1_awready),
        .o_awaddr     (slv1_awaddr),
        .o_awlen      (slv1_awlen),
        .o_awsize     (slv1_awsize),
        .o_awburst    (slv1_awburst),
        .o_awlock     (slv1_awlock),
        .o_awid       (slv1_awid),
        .o_wvalid     (slv1_wvalid),
        .o_wready     (slv1_wready),
        .o_wlast      (slv1_wlast),
        .o_wid        (slv1_wid),
        .o_wdata      (slv1_wdata),
        .o_wstrb      (slv1_wstrb),
        .o_bvalid     (slv1_bvalid),
        .o_bready     (slv1_bready),
        .o_bid        (slv1_bid),
        .o_bresp      (slv1_bresp),
        .o_arvalid    (slv1_arvalid),
        .o_arready    (slv1_arready),
        .o_araddr     (slv1_araddr),
        .o_arlen      (slv1_arlen),
        .o_arsize     (slv1_arsize),
        .o_arburst    (slv1_arburst),
        .o_arlock     (slv1_arlock),
        .o_arid       (slv1_arid),
        .o_rvalid     (slv1_rvalid),
        .o_rready     (slv1_rready),
        .o_rid        (slv1_rid),
        .o_rresp      (slv1_rresp),
        .o_rdata      (slv1_rdata),
        .o_rlast      (slv1_rlast)
    );

    ////////////////////////////////
    //slv2 interface
    ///////////////////////////////
    axi_crossbar_slv_if#(
        .AXI_ADDR_W       (AXI_ADDR_W),
        .AXI_ID_W         (AXI_ID_W),
        .AXI_DATA_W       (AXI_DATA_W),
        .BASE_ADDR        (SLV2_START_ADDR),
        .SLV_OSTDREQ_NUM  (SLV2_OSTDREQ_NUM),
        .SLV_OSTDREQ_SIZE (SLV2_OSTDREQ_SIZE),
        .AWCH_W           (AWCH_W),
        .WCH_W            (WCH_W),
        .BCH_W            (BCH_W),
        .ARCH_W           (ARCH_W),
        .RCH_W            (RCH_W)
    )
    slv2_if(
         //interface from switch
        .i_aclk       (aclk),
        .i_aresetn    (aresetn),
        .i_srst       (srst),
        .i_awvalid    (o_awvalid[2]),
        .i_awready    (o_awready[2]),
        .i_awch       (o_awch[2*AWCH_W+:AWCH_W]),
        .i_wvalid     (o_wvalid[2]),
        .i_wready     (o_wready[2]),
        .i_wlast      (o_wlast[2]),
        .i_wch        (o_wch[2*WCH_W+:WCH_W]),
        .i_bvalid     (o_bvalid[2]),
        .i_bready     (o_bready[2]),
        .i_bch        (o_bch[2*BCH_W+:BCH_W]),
        .i_arvalid    (o_arvalid[2]),
        .i_arready    (o_arready[2]),
        .i_arch       (o_arch[2*ARCH_W+:ARCH_W]),
        .i_rvalid     (o_rvalid[2]),
        .i_rready     (o_rready[2]),
        .i_rlast      (o_rlast[2]),
        .i_rch        (o_rch[2*RCH_W+:RCH_W]),
        //interface to slave
        .o_aclk       (slv2_aclk),
        .o_aresetn    (slv2_aresetn),
        .o_srst       (slv2_srst),
        .o_awvalid    (slv2_awvalid),
        .o_awready    (slv2_awready),
        .o_awaddr     (slv2_awaddr),
        .o_awlen      (slv2_awlen),
        .o_awsize     (slv2_awsize),
        .o_awburst    (slv2_awburst),
        .o_awlock     (slv2_awlock),
        .o_awid       (slv2_awid),
        .o_wvalid     (slv2_wvalid),
        .o_wready     (slv2_wready),
        .o_wlast      (slv2_wlast),
        .o_wid        (slv2_wid),
        .o_wdata      (slv2_wdata),
        .o_wstrb      (slv2_wstrb),
        .o_bvalid     (slv2_bvalid),
        .o_bready     (slv2_bready),
        .o_bid        (slv2_bid),
        .o_bresp      (slv2_bresp),
        .o_arvalid    (slv2_arvalid),
        .o_arready    (slv2_arready),
        .o_araddr     (slv2_araddr),
        .o_arlen      (slv2_arlen),
        .o_arsize     (slv2_arsize),
        .o_arburst    (slv2_arburst),
        .o_arlock     (slv2_arlock),
        .o_arid       (slv2_arid),
        .o_rvalid     (slv2_rvalid),
        .o_rready     (slv2_rready),
        .o_rid        (slv2_rid),
        .o_rresp      (slv2_rresp),
        .o_rdata      (slv2_rdata),
        .o_rlast      (slv2_rlast)
    );        



endmodule


`resetall